.title KiCad schematic
R1 NODE1 NODE2 1k
V1 NODE1 0 1
R2 NODE2 0 2k
.control
    op
    print v(node2)
.endc
.end
